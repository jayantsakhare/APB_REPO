class apb_configuration;
endclass
